module main

import os
import json
import term
import rand

const json_string = '[{"name":"Aatrox","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2013,"species":"Darkin","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Aatrox.png","gender":"Male","resource":"Blood Well"},{"name":"Ahri","roles":["Assassin","Mage"],"lanes":["Middle"],"release_date":2011,"species":"Vastayan","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ahri.png","gender":"Female","resource":"Mana"},{"name":"Akali","roles":["Assassin"],"lanes":["Middle","Top"],"release_date":2010,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Akali.png","gender":"Female","resource":"Energy"},{"name":"Akshan","roles":["Assassin","Marksman"],"lanes":["Middle"],"release_date":2021,"species":"Human","region":"Shurima","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Akshan.png","gender":"Male","resource":"Mana"},{"name":"Alistar","roles":["Tank","Support"],"lanes":["Support"],"release_date":2009,"species":"Minotaur","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Alistar.png","gender":"Male","resource":"Mana"},{"name":"Amumu","roles":["Tank","Mage"],"lanes":["Support"],"release_date":2009,"species":"Unknown","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Amumu.png","gender":"Unknown","resource":"Mana"},{"name":"Anivia","roles":["Mage","Support"],"lanes":["Middle"],"release_date":2009,"species":"Spirit God","region":"Freljord","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Anivia.png","gender":"Female","resource":"Mana"},{"name":"Annie","roles":["Mage"],"lanes":["Middle"],"release_date":2009,"species":"Human","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Annie.png","gender":"Female","resource":"Mana"},{"name":"Aphelios","roles":["Marksman"],"lanes":["Bottom"],"release_date":2019,"species":"Human","region":"Targon","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Aphelios.png","gender":"Male","resource":"Mana"},{"name":"Ashe","roles":["Marksman","Support"],"lanes":["Support","Bottom"],"release_date":2009,"species":"Human","region":"Freljord","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ashe.png","gender":"Female","resource":"Mana"},{"name":"Aurelion Sol","roles":["Mage"],"lanes":["Middle"],"release_date":2016,"species":"Celestial","region":"Targon","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/AurelionSol.png","gender":"Male","resource":"Mana"},{"name":"Azir","roles":["Mage","Marksman"],"lanes":["Middle"],"release_date":2014,"species":"God-Warrior","region":"Shurima","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Azir.png","gender":"Male","resource":"Mana"},{"name":"Bard","roles":["Mage","Support"],"lanes":["Support"],"release_date":2015,"species":"Celestial","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Bard.png","gender":"Male","resource":"Mana"},{"name":"Bel\'Veth","roles":["Fighter"],"lanes":["Jungle"],"release_date":2022,"species":"Voidborn","region":"Void","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.11.1/img/champion/Belveth.png","gender":"Unknown","resource":"Mana"},{"name":"Blitzcrank","roles":["Fighter","Tank"],"lanes":["Support"],"release_date":2009,"species":"Golem","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Blitzcrank.png","gender":"Unknown","resource":"Mana"},{"name":"Brand","roles":["Mage"],"lanes":["Support"],"release_date":2011,"species":"Human","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Brand.png","gender":"Male","resource":"Mana"},{"name":"Braum","roles":["Tank","Support"],"lanes":["Support"],"release_date":2014,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Braum.png","gender":"Male","resource":"Mana"},{"name":"Caitlyn","roles":["Marksman"],"lanes":["Bottom"],"release_date":2011,"species":"Human","region":"Piltover","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Caitlyn.png","gender":"Female","resource":"Mana"},{"name":"Camille","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2016,"species":"Human","region":"Piltover","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Camille.png","gender":"Female","resource":"Mana"},{"name":"Cassiopeia","roles":["Mage"],"lanes":["Middle"],"release_date":2010,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Cassiopeia.png","gender":"Female","resource":"Mana"},{"name":"Cho\'Gath","roles":["Tank","Mage"],"lanes":["Top"],"release_date":2009,"species":"Voidborn","region":"Void","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Chogath.png","gender":"Male","resource":"Mana"},{"name":"Corki","roles":["Marksman"],"lanes":["Middle"],"release_date":2009,"species":"Yordle","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Corki.png","gender":"Male","resource":"Mana"},{"name":"Darius","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2012,"species":"Human","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Darius.png","gender":"Male","resource":"Mana"},{"name":"Diana","roles":["Fighter","Mage"],"lanes":["Jungle"],"release_date":2012,"species":"Aspect Host","region":"Targon","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Diana.png","gender":"Female","resource":"Mana"},{"name":"Dr. Mundo","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2009,"species":"Human","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/DrMundo.png","gender":"Male","resource":"Health"},{"name":"Draven","roles":["Marksman"],"lanes":["Bottom"],"release_date":2012,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Draven.png","gender":"Male","resource":"Mana"},{"name":"Ekko","roles":["Fighter","Assassin"],"lanes":["Jungle","Middle"],"release_date":2015,"species":"Human","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ekko.png","gender":"Male","resource":"Mana"},{"name":"Elise","roles":["Fighter","Mage"],"lanes":["Jungle"],"release_date":2012,"species":"Human","region":"Shadow Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Elise.png","gender":"Female","resource":"Mana"},{"name":"Evelynn","roles":["Assassin","Mage"],"lanes":["Jungle"],"release_date":2009,"species":"Demon","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Evelynn.png","gender":"Female","resource":"Mana"},{"name":"Ezreal","roles":["Mage","Marksman"],"lanes":["Bottom"],"release_date":2010,"species":"Human","region":"Piltover","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ezreal.png","gender":"Male","resource":"Mana"},{"name":"Fiddlesticks","roles":["Mage","Support"],"lanes":["Jungle"],"release_date":2009,"species":"Demon","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Fiddlesticks.png","gender":"Unknown","resource":"Mana"},{"name":"Fiora","roles":["Fighter","Assassin"],"lanes":["Top"],"release_date":2012,"species":"Human","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Fiora.png","gender":"Female","resource":"Mana"},{"name":"Fizz","roles":["Fighter","Assassin"],"lanes":["Middle"],"release_date":2011,"species":"Yordle","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Fizz.png","gender":"Male","resource":"Mana"},{"name":"Galio","roles":["Tank","Mage"],"lanes":["Middle"],"release_date":2010,"species":"Golem","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Galio.png","gender":"Unknown","resource":"Mana"},{"name":"Gangplank","roles":["Fighter"],"lanes":["Top"],"release_date":2009,"species":"Human","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Gangplank.png","gender":"Male","resource":"Mana"},{"name":"Garen","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2010,"species":"Human","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Garen.png","gender":"Male","resource":"None"},{"name":"Gnar","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2014,"species":"Yordle","region":"Freljord","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Gnar.png","gender":"Male","resource":"Rage"},{"name":"Gragas","roles":["Fighter","Mage"],"lanes":["Top"],"release_date":2010,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Gragas.png","gender":"Male","resource":"Mana"},{"name":"Graves","roles":["Marksman"],"lanes":["Jungle"],"release_date":2011,"species":"Human","region":"Bilgewater","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Graves.png","gender":"Male","resource":"Mana"},{"name":"Gwen","roles":["Fighter","Assassin"],"lanes":["Top"],"release_date":2021,"species":"Human","region":"Shadow Isles","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Gwen.png","gender":"Female","resource":"Mana"},{"name":"Hecarim","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2012,"species":"Wraith","region":"Shadow Isles","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Hecarim.png","gender":"Male","resource":"Mana"},{"name":"Heimerdinger","roles":["Mage","Support"],"lanes":["Support"],"release_date":2009,"species":"Yordle","region":"Piltover","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Heimerdinger.png","gender":"Male","resource":"Mana"},{"name":"Illaoi","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2015,"species":"Human","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Illaoi.png","gender":"Female","resource":"Mana"},{"name":"Irelia","roles":["Fighter","Assassin"],"lanes":["Middle","Top"],"release_date":2010,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Irelia.png","gender":"Female","resource":"Mana"},{"name":"Ivern","roles":["Mage","Support"],"lanes":["Jungle"],"release_date":2016,"species":"Human","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ivern.png","gender":"Male","resource":"Mana"},{"name":"Janna","roles":["Mage","Support"],"lanes":["Support"],"release_date":2009,"species":"Spirit God","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Janna.png","gender":"Female","resource":"Mana"},{"name":"Jarvan IV","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2011,"species":"Human","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/JarvanIV.png","gender":"Male","resource":"Mana"},{"name":"Jax","roles":["Fighter","Assassin"],"lanes":["Top"],"release_date":2009,"species":"Unknown","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Jax.png","gender":"Unknown","resource":"Mana"},{"name":"Jayce","roles":["Fighter","Marksman"],"lanes":["Top"],"release_date":2012,"species":"Human","region":"Piltover","range_type":["Melee","Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Jayce.png","gender":"Male","resource":"Mana"},{"name":"Jhin","roles":["Mage","Marksman"],"lanes":["Bottom"],"release_date":2016,"species":"Human","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Jhin.png","gender":"Male","resource":"Mana"},{"name":"Jinx","roles":["Marksman"],"lanes":["Bottom"],"release_date":2013,"species":"Human","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Jinx.png","gender":"Female","resource":"Mana"},{"name":"K\'Sante","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2022,"species":"Human","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.21.1/img/champion/KSante.png","gender":"Male","resource":"Mana"},{"name":"Kai\'Sa","roles":["Marksman"],"lanes":["Bottom"],"release_date":2018,"species":"Human","region":"Void","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kaisa.png","gender":"Female","resource":"Mana"},{"name":"Kalista","roles":["Marksman"],"lanes":["Bottom"],"release_date":2014,"species":"Wraith","region":"Shadow Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kalista.png","gender":"Female","resource":"Mana"},{"name":"Karma","roles":["Mage","Support"],"lanes":["Support"],"release_date":2011,"species":"Human","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Karma.png","gender":"Female","resource":"Mana"},{"name":"Karthus","roles":["Mage"],"lanes":["Jungle"],"release_date":2009,"species":"Wraith","region":"Shadow Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Karthus.png","gender":"Male","resource":"Mana"},{"name":"Kassadin","roles":["Assassin","Mage"],"lanes":["Middle"],"release_date":2009,"species":"Human","region":"Void","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kassadin.png","gender":"Male","resource":"Mana"},{"name":"Katarina","roles":["Assassin","Mage"],"lanes":["Middle"],"release_date":2009,"species":"Human","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Katarina.png","gender":"Female","resource":"None"},{"name":"Kayle","roles":["Fighter","Support"],"lanes":["Top"],"release_date":2009,"species":"Human","region":"Targon","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kayle.png","gender":"Female","resource":"Mana"},{"name":"Kayn","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2017,"species":"Darkin","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kayn.png","gender":"Male","resource":"Mana"},{"name":"Kennen","roles":["Mage","Marksman"],"lanes":["Top"],"release_date":2010,"species":"Yordle","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kennen.png","gender":"Male","resource":"Energy"},{"name":"Kha\'Zix","roles":["Assassin"],"lanes":["Jungle"],"release_date":2012,"species":"Voidborn","region":"Void","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Khazix.png","gender":"Male","resource":"Mana"},{"name":"Kindred","roles":["Marksman"],"lanes":["Jungle"],"release_date":2015,"species":"Spirit God","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kindred.png","gender":"Unknown","resource":"Mana"},{"name":"Kled","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2016,"species":"Yordle","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Kled.png","gender":"Male","resource":"Courage"},{"name":"Kog\'Maw","roles":["Mage","Marksman"],"lanes":["Bottom"],"release_date":2010,"species":"Voidborn","region":"Void","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/KogMaw.png","gender":"Male","resource":"Mana"},{"name":"LeBlanc","roles":["Assassin","Mage"],"lanes":["Middle"],"release_date":2010,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Leblanc.png","gender":"Female","resource":"Mana"},{"name":"Lee Sin","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2011,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/LeeSin.png","gender":"Male","resource":"Energy"},{"name":"Leona","roles":["Tank","Support"],"lanes":["Support"],"release_date":2011,"species":"Aspect Host","region":"Targon","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Leona.png","gender":"Female","resource":"Mana"},{"name":"Lillia","roles":["Fighter","Mage"],"lanes":["Jungle"],"release_date":2020,"species":"Spirit","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Lillia.png","gender":"Female","resource":"Mana"},{"name":"Lissandra","roles":["Mage"],"lanes":["Middle"],"release_date":2013,"species":"Human","region":"Freljord","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Lissandra.png","gender":"Female","resource":"Mana"},{"name":"Lucian","roles":["Marksman"],"lanes":["Bottom"],"release_date":2013,"species":"Human","region":"Blessed Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Lucian.png","gender":"Male","resource":"Mana"},{"name":"Lulu","roles":["Mage","Support"],"lanes":["Support"],"release_date":2012,"species":"Yordle","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Lulu.png","gender":"Female","resource":"Mana"},{"name":"Lux","roles":["Mage","Support"],"lanes":["Support","Middle"],"release_date":2010,"species":"Human","region":"Demacia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Lux.png","gender":"Female","resource":"Mana"},{"name":"Malphite","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2009,"species":"Golem","region":"Ixtal","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Malphite.png","gender":"Male","resource":"Mana"},{"name":"Malzahar","roles":["Assassin","Mage"],"lanes":["Middle"],"release_date":2010,"species":"Human","region":"Void","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Malzahar.png","gender":"Male","resource":"Mana"},{"name":"Maokai","roles":["Tank","Mage"],"lanes":["Support"],"release_date":2011,"species":"Spirit","region":"Shadow Isles","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Maokai.png","gender":"Unknown","resource":"Mana"},{"name":"Master Yi","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2009,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/MasterYi.png","gender":"Male","resource":"Mana"},{"name":"Miss Fortune","roles":["Marksman"],"lanes":["Bottom"],"release_date":2010,"species":"Human","region":"Bilgewater","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/MissFortune.png","gender":"Female","resource":"Mana"},{"name":"Mordekaiser","roles":["Fighter"],"lanes":["Jungle","Top"],"release_date":2010,"species":"Revenant","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Mordekaiser.png","gender":"Male","resource":"Shield"},{"name":"Morgana","roles":["Mage","Support"],"lanes":["Support"],"release_date":2009,"species":"Human","region":"Targon","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Morgana.png","gender":"Female","resource":"Mana"},{"name":"Nami","roles":["Mage","Support"],"lanes":["Support"],"release_date":2012,"species":"Vastayan","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nami.png","gender":"Female","resource":"Mana"},{"name":"Nasus","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2009,"species":"God-Warrior","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nasus.png","gender":"Male","resource":"Mana"},{"name":"Nautilus","roles":["Fighter","Tank"],"lanes":["Support"],"release_date":2012,"species":"Revenant","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nautilus.png","gender":"Male","resource":"Mana"},{"name":"Neeko","roles":["Mage","Support"],"lanes":["Middle"],"release_date":2018,"species":"Vastayan","region":"Ixtal","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Neeko.png","gender":"Female","resource":"Mana"},{"name":"Nidalee","roles":["Assassin","Mage"],"lanes":["Jungle"],"release_date":2009,"species":"Human","region":"Ixtal","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nidalee.png","gender":"Female","resource":"Mana"},{"name":"Nilah","roles":["Fighter","Assassin"],"lanes":["Bottom"],"release_date":2022,"species":"Human","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.13.1/img/champion/Nilah.png","gender":"Female","resource":"Mana"},{"name":"Nocturne","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2011,"species":"Demon","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nocturne.png","gender":"Unknown","resource":"Mana"},{"name":"Nunu & Willump","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2009,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Nunu.png","gender":"Male","resource":"Mana"},{"name":"Olaf","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2010,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Olaf.png","gender":"Male","resource":"Mana"},{"name":"Orianna","roles":["Mage","Support"],"lanes":["Middle"],"release_date":2011,"species":"Golem","region":"Piltover","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Orianna.png","gender":"Female","resource":"Mana"},{"name":"Ornn","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2017,"species":"Spirit God","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ornn.png","gender":"Male","resource":"Mana"},{"name":"Pantheon","roles":["Fighter","Assassin"],"lanes":["Support"],"release_date":2010,"species":"Aspect Host","region":"Targon","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Pantheon.png","gender":"Male","resource":"Mana"},{"name":"Poppy","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2010,"species":"Yordle","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Poppy.png","gender":"Female","resource":"Mana"},{"name":"Pyke","roles":["Assassin","Support"],"lanes":["Support"],"release_date":2018,"species":"Revenant","region":"Bilgewater","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Pyke.png","gender":"Male","resource":"Mana"},{"name":"Qiyana","roles":["Fighter","Assassin"],"lanes":["Middle"],"release_date":2019,"species":"Human","region":"Ixtal","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Qiyana.png","gender":"Female","resource":"Mana"},{"name":"Quinn","roles":["Assassin","Marksman"],"lanes":["Top"],"release_date":2013,"species":"Human","region":"Demacia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Quinn.png","gender":"Female","resource":"Mana"},{"name":"Rakan","roles":["Support"],"lanes":["Support"],"release_date":2017,"species":"Vastayan","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Rakan.png","gender":"Male","resource":"Mana"},{"name":"Rammus","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2009,"species":"Unknown","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Rammus.png","gender":"Male","resource":"Mana"},{"name":"Rek\'Sai","roles":["Fighter"],"lanes":["Jungle"],"release_date":2014,"species":"Voidborn","region":"Void","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/RekSai.png","gender":"Female","resource":"Rage"},{"name":"Rell","roles":["Tank"],"lanes":["Support"],"release_date":2020,"species":"Human","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Rell.png","gender":"Female","resource":"Mana"},{"name":"Renata Glasc","roles":["Mage","Support"],"lanes":["Support"],"release_date":2022,"species":"Human","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.7.1/img/champion/Renata.png","gender":"Female","resource":"Mana"},{"name":"Renekton","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2011,"species":"God-Warrior","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Renekton.png","gender":"Male","resource":"Fury"},{"name":"Rengar","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2012,"species":"Vastayan","region":"Ixtal","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Rengar.png","gender":"Male","resource":"Ferocity"},{"name":"Riven","roles":["Fighter","Assassin"],"lanes":["Top"],"release_date":2011,"species":"Human","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Riven.png","gender":"Female","resource":"None"},{"name":"Rumble","roles":["Fighter","Mage"],"lanes":["Middle","Top"],"release_date":2011,"species":"Yordle","region":"Bandle City","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Rumble.png","gender":"Male","resource":"Heat"},{"name":"Ryze","roles":["Fighter","Mage"],"lanes":["Middle"],"release_date":2009,"species":"Human","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ryze.png","gender":"Male","resource":"Mana"},{"name":"Samira","roles":["Marksman"],"lanes":["Bottom"],"release_date":2020,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Samira.png","gender":"Female","resource":"Mana"},{"name":"Sejuani","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2012,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sejuani.png","gender":"Female","resource":"Mana"},{"name":"Senna","roles":["Marksman","Support"],"lanes":["Support"],"release_date":2019,"species":"Human","region":"Blessed Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Senna.png","gender":"Female","resource":"Mana"},{"name":"Seraphine","roles":["Mage","Support"],"lanes":["Support"],"release_date":2020,"species":"Human","region":"Piltover","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Seraphine.png","gender":"Female","resource":"Mana"},{"name":"Sett","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2020,"species":"Vastayan","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sett.png","gender":"Male","resource":"Grit"},{"name":"Shaco","roles":["Assassin"],"lanes":["Jungle"],"release_date":2009,"species":"Spirit","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Shaco.png","gender":"Male","resource":"Mana"},{"name":"Shen","roles":["Tank"],"lanes":["Top"],"release_date":2010,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Shen.png","gender":"Male","resource":"Energy"},{"name":"Shyvana","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2011,"species":"Terrestrial Dragon","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Shyvana.png","gender":"Female","resource":"Fury"},{"name":"Singed","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2009,"species":"Human","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Singed.png","gender":"Male","resource":"Mana"},{"name":"Sion","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2009,"species":"Revenant","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sion.png","gender":"Male","resource":"Mana"},{"name":"Sivir","roles":["Marksman"],"lanes":["Bottom"],"release_date":2009,"species":"Human","region":"Shurima","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sivir.png","gender":"Female","resource":"Mana"},{"name":"Skarner","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2011,"species":"Brackern","region":"Shurima","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Skarner.png","gender":"Male","resource":"Mana"},{"name":"Sona","roles":["Mage","Support"],"lanes":["Support"],"release_date":2010,"species":"Human","region":"Demacia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sona.png","gender":"Female","resource":"Mana"},{"name":"Soraka","roles":["Mage","Support"],"lanes":["Support"],"release_date":2009,"species":"Celestial","region":"Targon","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Soraka.png","gender":"Female","resource":"Mana"},{"name":"Swain","roles":["Fighter","Mage"],"lanes":["Support","Middle"],"release_date":2010,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Swain.png","gender":"Male","resource":"Mana"},{"name":"Sylas","roles":["Assassin","Mage"],"lanes":["Jungle","Middle"],"release_date":2019,"species":"Human","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Sylas.png","gender":"Male","resource":"Mana"},{"name":"Syndra","roles":["Mage","Support"],"lanes":["Middle"],"release_date":2012,"species":"Human","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Syndra.png","gender":"Female","resource":"Mana"},{"name":"Tahm Kench","roles":["Tank","Support"],"lanes":["Top"],"release_date":2015,"species":"Demon","region":"Runeterra","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/TahmKench.png","gender":"Male","resource":"Mana"},{"name":"Taliyah","roles":["Mage","Support"],"lanes":["Jungle","Middle"],"release_date":2016,"species":"Human","region":"Shurima","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Taliyah.png","gender":"Female","resource":"Mana"},{"name":"Talon","roles":["Assassin"],"lanes":["Middle"],"release_date":2011,"species":"Human","region":"Noxus","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Talon.png","gender":"Male","resource":"Mana"},{"name":"Taric","roles":["Fighter","Support"],"lanes":["Support"],"release_date":2009,"species":"Aspect Host","region":"Targon","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Taric.png","gender":"Male","resource":"Mana"},{"name":"Teemo","roles":["Assassin","Marksman"],"lanes":["Top"],"release_date":2009,"species":"Yordle","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Teemo.png","gender":"Male","resource":"Mana"},{"name":"Thresh","roles":["Fighter","Support"],"lanes":["Support"],"release_date":2013,"species":"Wraith","region":"Shadow Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Thresh.png","gender":"Male","resource":"Mana"},{"name":"Tristana","roles":["Assassin","Marksman"],"lanes":["Bottom"],"release_date":2009,"species":"Yordle","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Tristana.png","gender":"Female","resource":"Mana"},{"name":"Trundle","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2010,"species":"Troll","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Trundle.png","gender":"Male","resource":"Mana"},{"name":"Tryndamere","roles":["Fighter","Assassin"],"lanes":["Top"],"release_date":2009,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Tryndamere.png","gender":"Male","resource":"Fury"},{"name":"Twisted Fate","roles":["Mage"],"lanes":["Middle"],"release_date":2009,"species":"Human","region":"Bilgewater","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/TwistedFate.png","gender":"Male","resource":"Mana"},{"name":"Twitch","roles":["Assassin","Marksman"],"lanes":["Bottom"],"release_date":2009,"species":"Plague Rat","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Twitch.png","gender":"Male","resource":"Mana"},{"name":"Udyr","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2009,"species":"Human","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.17.1/img/champion/Udyr.png","gender":"Male","resource":"Mana"},{"name":"Urgot","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2010,"species":"Human","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Urgot.png","gender":"Male","resource":"Mana"},{"name":"Varus","roles":["Mage","Marksman"],"lanes":["Middle","Bottom"],"release_date":2012,"species":"Darkin","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Varus.png","gender":"Male","resource":"Mana"},{"name":"Vayne","roles":["Assassin","Marksman"],"lanes":["Bottom"],"release_date":2011,"species":"Human","region":"Demacia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Vayne.png","gender":"Female","resource":"Mana"},{"name":"Veigar","roles":["Mage"],"lanes":["Middle"],"release_date":2009,"species":"Yordle","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Veigar.png","gender":"Male","resource":"Mana"},{"name":"Vel\'Koz","roles":["Mage"],"lanes":["Support"],"release_date":2014,"species":"Voidborn","region":"Void","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Velkoz.png","gender":"Male","resource":"Mana"},{"name":"Vex","roles":["Mage"],"lanes":["Middle"],"release_date":2021,"species":"Yordle","region":"Shadow Isles","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Vex.png","gender":"Female","resource":"Mana"},{"name":"Vi","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2012,"species":"Human","region":"Piltover","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Vi.png","gender":"Female","resource":"Mana"},{"name":"Viego","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2021,"species":"Wraith","region":"Shadow Isles","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Viego.png","gender":"Male","resource":"None"},{"name":"Viktor","roles":["Mage"],"lanes":["Middle"],"release_date":2011,"species":"Human","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Viktor.png","gender":"Male","resource":"Mana"},{"name":"Vladimir","roles":["Mage"],"lanes":["Middle"],"release_date":2010,"species":"Human","region":"Noxus","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Vladimir.png","gender":"Male","resource":"Crimson Rush"},{"name":"Volibear","roles":["Fighter","Tank"],"lanes":["Jungle","Top"],"release_date":2011,"species":"Spirit God","region":"Freljord","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Volibear.png","gender":"Male","resource":"Mana"},{"name":"Warwick","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2009,"species":"Human","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Warwick.png","gender":"Male","resource":"Mana"},{"name":"Wukong","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2011,"species":"Vastayan","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/MonkeyKing.png","gender":"Male","resource":"Mana"},{"name":"Xayah","roles":["Marksman"],"lanes":["Bottom"],"release_date":2017,"species":"Vastayan","region":"Ionia","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Xayah.png","gender":"Female","resource":"Mana"},{"name":"Xerath","roles":["Mage"],"lanes":["Support"],"release_date":2011,"species":"Baccai","region":"Shurima","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Xerath.png","gender":"Male","resource":"Mana"},{"name":"Xin Zhao","roles":["Fighter","Assassin"],"lanes":["Jungle"],"release_date":2010,"species":"Human","region":"Demacia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/XinZhao.png","gender":"Male","resource":"Mana"},{"name":"Yasuo","roles":["Fighter","Assassin"],"lanes":["Middle","Top"],"release_date":2013,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Yasuo.png","gender":"Male","resource":"Flow"},{"name":"Yone","roles":["Fighter","Assassin"],"lanes":["Middle","Top"],"release_date":2020,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Yone.png","gender":"Male","resource":"Flow"},{"name":"Yorick","roles":["Fighter","Tank"],"lanes":["Top"],"release_date":2011,"species":"Human","region":"Shadow Isles","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Yorick.png","gender":"Male","resource":"Mana"},{"name":"Yuumi","roles":["Mage","Support"],"lanes":["Support"],"release_date":2019,"species":"Cat","region":"Bandle City","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Yuumi.png","gender":"Female","resource":"Mana"},{"name":"Zac","roles":["Fighter","Tank"],"lanes":["Jungle"],"release_date":2013,"species":"Golem","region":"Zaun","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Zac.png","gender":"Male","resource":"Health"},{"name":"Zed","roles":["Assassin"],"lanes":["Jungle","Middle"],"release_date":2012,"species":"Human","region":"Ionia","range_type":["Melee"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Zed.png","gender":"Male","resource":"Energy"},{"name":"Zeri","roles":["Marksman"],"lanes":["Bottom"],"release_date":2022,"species":"Human","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/12.7.1/img/champion/Zeri.png","gender":"Female","resource":"Mana"},{"name":"Ziggs","roles":["Mage"],"lanes":["Middle"],"release_date":2012,"species":"Yordle","region":"Zaun","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Ziggs.png","gender":"Male","resource":"Mana"},{"name":"Zilean","roles":["Mage","Support"],"lanes":["Support"],"release_date":2009,"species":"Human","region":"Runeterra","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Zilean.png","gender":"Male","resource":"Mana"},{"name":"Zoe","roles":["Mage","Support"],"lanes":["Middle"],"release_date":2017,"species":"Aspect Host","region":"Targon","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Zoe.png","gender":"Female","resource":"Mana"},{"name":"Zyra","roles":["Mage","Support"],"lanes":["Support"],"release_date":2012,"species":"Unknown","region":"Ixtal","range_type":["Ranged"],"portrait":"https://ddragon.leagueoflegends.com/cdn/11.23.1/img/champion/Zyra.png","gender":"Female","resource":"Mana"}]'

struct Champion {
	name         string
	roles        []string
	lanes        []string
	release_date int
	species      string
	region       string
	range_type   []string
	portrait     string
	gender       string
	resource     string
}

const green = '\033[92m'

const yellow = '\033[93m'

const red = '\033[91m'

const end = '\033[0m'

const blue = '\033[94m'

enum GuessResult {
	registered
	already_guessed
	success
	not_found
}

struct App {
	all_champs []Champion
mut:
	to_guess Champion
	guesses  []Champion
}

fn main() {
	all_champs := load_champs()
	mut app := &App{
		all_champs: all_champs
		to_guess: rand.choose[Champion](all_champs, 1)![0]
	}

	println('Start by guessing a champion name.')
	mut guess_count := 0
	for {
		input := os.input('(${guess_count}) Your guess: ')
		result := app.guess(input)

		if input.to_lower() == 'end' {
			println('The Champion was ${app.to_guess.name}.')
			break
		}

		match result {
			.registered {
				guess_count += 1
				app.print_guessed()
			}
			.success {
				app.print_guessed()
				x, _ := term.get_terminal_size()
				println('')
				println(term.yellow('${' '.repeat((x - 9) / 2)}Congrats!'))
				println(term.yellow('${' '.repeat((x - 18 - (guess_count + 1).str().len) / 2)}It took you ${
					guess_count + 1} guesses.'))
				println('')
				break
			}
			else {
				println('Try again!')
			}
		}
	}
}

fn (a App) print_guessed() {
	term.clear()

	pr(blue, 'Name')
	pr(blue, 'Gender')
	pr(blue, 'Lanes')
	pr(blue, 'Species')
	pr(blue, 'Resource')
	pr(blue, 'Range Type')
	pr(blue, 'Region')
	pr(blue, 'Release')
	println('')

	for c in a.guesses {
		pr(blue, c.name)
		pr_sgl(c.gender, a.to_guess.gender)
		pr_arr(c.lanes, a.to_guess.lanes)
		pr_sgl(c.species, a.to_guess.species)
		pr_sgl(c.resource, a.to_guess.resource)
		pr_arr(c.range_type, a.to_guess.range_type)
		pr_sgl(c.region, a.to_guess.region)

		if c.release_date == a.to_guess.release_date {
			pr(green, '${c.release_date}')
		} else {
			if c.release_date > a.to_guess.release_date {
				pr(red, '${c.release_date} 🔽')
			} else {
				pr(red, '${c.release_date} 🔼')
			}
		}
		println('')
	}
}

fn pr_sgl(a string, b string) {
	if a == b {
		pr(green, a)
	} else {
		pr(red, a)
	}
}

fn pr(color string, field string) {
	print('${color}${field:-16}${end}')
}

fn pr_arr(guess []string, a []string) {
	if a == guess {
		pr(green, guess.join(', '))
	} else {
		if guess.any(it in a) {
			pr(yellow, guess.join(', '))
		} else {
			pr(red, guess.join(', '))
		}
	}
}

fn (mut a App) guess(input string) GuessResult {
	champ := a.find_champ(input) or { return .not_found }

	if a.to_guess.name == champ.name {
		a.guesses << champ
		return .success
	} else if champ in a.guesses {
		return .already_guessed
	}

	a.guesses << champ
	return .registered
}

fn (a App) find_champ(name string) !Champion {
	for i in a.all_champs {
		if i.name.to_lower().starts_with(name.to_lower()) {
			return i
		}
	}
	return error('No champion found')
}

fn load_champs() []Champion {
	champs := json.decode([]Champion, json_string) or { [] }
	return champs
}
